-- XXX
-- Aaka Fosfor, 2020
-- https://github.com/AakaFosfor/hdl_cores
--
-- state: draft

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity XXX is
  generic (
    G_CLK_FREQUENCY : real; -- in Hz
    XXX
  );
  port (
    Clk_ik   : in  std_logic;
    Reset_ir : in  std_logic;
    XXX
  );
end entity;

architecture RTL of XXX is

  XXX

begin

  XXX

end architecture;
